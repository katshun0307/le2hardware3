library verilog;
use verilog.vl_types.all;
entity main_vlg_tst is
end main_vlg_tst;
