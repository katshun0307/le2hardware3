library verilog;
use verilog.vl_types.all;
entity xor1616_vlg_tst is
end xor1616_vlg_tst;
