library verilog;
use verilog.vl_types.all;
entity sub16_vlg_tst is
end sub16_vlg_tst;
